// top level module for project
// literally nothing yet

module tic_tac_toe()
endmodule
