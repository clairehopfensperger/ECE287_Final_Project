// completely empty module, created to acknowledge that we want a display module

module display();

endmodule
